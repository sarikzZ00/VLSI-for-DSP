module cosine_LUT (
    input [7:0] phase,
    output logic signed [7:0] cosine_value
);

    always_comb begin
        case (phase)
            8'd0: cosine_value = 127;
            8'd1: cosine_value = 127;
            8'd2: cosine_value = 127;
            8'd3: cosine_value = 127;
            8'd4: cosine_value = 127;
            8'd5: cosine_value = 127;
            8'd6: cosine_value = 127;
            8'd7: cosine_value = 126;
            8'd8: cosine_value = 126;
            8'd9: cosine_value = 125;
            8'd10: cosine_value = 124;
            8'd11: cosine_value = 123;
            8'd12: cosine_value = 122;
            8'd13: cosine_value = 122;
            8'd14: cosine_value = 121;
            8'd15: cosine_value = 119;
            8'd16: cosine_value = 118;
            8'd17: cosine_value = 117;
            8'd18: cosine_value = 116;
            8'd19: cosine_value = 114;
            8'd20: cosine_value = 113;
            8'd21: cosine_value = 111;
            8'd22: cosine_value = 110;
            8'd23: cosine_value = 108;
            8'd24: cosine_value = 106;
            8'd25: cosine_value = 105;
            8'd26: cosine_value = 103;
            8'd27: cosine_value = 101;
            8'd28: cosine_value = 99;
            8'd29: cosine_value = 97;
            8'd30: cosine_value = 95;
            8'd31: cosine_value = 93;
            8'd32: cosine_value = 91;
            8'd33: cosine_value = 88;
            8'd34: cosine_value = 86;
            8'd35: cosine_value = 84;
            8'd36: cosine_value = 81;
            8'd37: cosine_value = 79;
            8'd38: cosine_value = 76;
            8'd39: cosine_value = 74;
            8'd40: cosine_value = 71;
            8'd41: cosine_value = 68;
            8'd42: cosine_value = 66;
            8'd43: cosine_value = 63;
            8'd44: cosine_value = 60;
            8'd45: cosine_value = 58;
            8'd46: cosine_value = 55;
            8'd47: cosine_value = 52;
            8'd48: cosine_value = 49;
            8'd49: cosine_value = 46;
            8'd50: cosine_value = 43;
            8'd51: cosine_value = 40;
            8'd52: cosine_value = 37;
            8'd53: cosine_value = 34;
            8'd54: cosine_value = 31;
            8'd55: cosine_value = 28;
            8'd56: cosine_value = 25;
            8'd57: cosine_value = 22;
            8'd58: cosine_value = 19;
            8'd59: cosine_value = 16;
            8'd60: cosine_value = 13;
            8'd61: cosine_value = 9;
            8'd62: cosine_value = 6;
            8'd63: cosine_value = 3;
            8'd64: cosine_value = 0;
            8'd65: cosine_value = -3;
            8'd66: cosine_value = -6;
            8'd67: cosine_value = -9;
            8'd68: cosine_value = -13;
            8'd69: cosine_value = -16;
            8'd70: cosine_value = -19;
            8'd71: cosine_value = -22;
            8'd72: cosine_value = -25;
            8'd73: cosine_value = -28;
            8'd74: cosine_value = -31;
            8'd75: cosine_value = -34;
            8'd76: cosine_value = -37;
            8'd77: cosine_value = -40;
            8'd78: cosine_value = -43;
            8'd79: cosine_value = -46;
            8'd80: cosine_value = -49;
            8'd81: cosine_value = -52;
            8'd82: cosine_value = -55;
            8'd83: cosine_value = -58;
            8'd84: cosine_value = -60;
            8'd85: cosine_value = -63;
            8'd86: cosine_value = -66;
            8'd87: cosine_value = -68;
            8'd88: cosine_value = -71;
            8'd89: cosine_value = -74;
            8'd90: cosine_value = -76;
            8'd91: cosine_value = -79;
            8'd92: cosine_value = -81;
            8'd93: cosine_value = -84;
            8'd94: cosine_value = -86;
            8'd95: cosine_value = -88;
            8'd96: cosine_value = -91;
            8'd97: cosine_value = -93;
            8'd98: cosine_value = -95;
            8'd99: cosine_value = -97;
            8'd100: cosine_value = -99;
            8'd101: cosine_value = -101;
            8'd102: cosine_value = -103;
            8'd103: cosine_value = -105;
            8'd104: cosine_value = -106;
            8'd105: cosine_value = -108;
            8'd106: cosine_value = -110;
            8'd107: cosine_value = -111;
            8'd108: cosine_value = -113;
            8'd109: cosine_value = -114;
            8'd110: cosine_value = -116;
            8'd111: cosine_value = -117;
            8'd112: cosine_value = -118;
            8'd113: cosine_value = -119;
            8'd114: cosine_value = -121;
            8'd115: cosine_value = -122;
            8'd116: cosine_value = -122;
            8'd117: cosine_value = -123;
            8'd118: cosine_value = -124;
            8'd119: cosine_value = -125;
            8'd120: cosine_value = -126;
            8'd121: cosine_value = -126;
            8'd122: cosine_value = -127;
            8'd123: cosine_value = -127;
            8'd124: cosine_value = -127;
            8'd125: cosine_value = -128;
            8'd126: cosine_value = -128;
            8'd127: cosine_value = -128;
            8'd128: cosine_value = -128;
            8'd129: cosine_value = -128;
            8'd130: cosine_value = -128;
            8'd131: cosine_value = -128;
            8'd132: cosine_value = -127;
            8'd133: cosine_value = -127;
            8'd134: cosine_value = -127;
            8'd135: cosine_value = -126;
            8'd136: cosine_value = -126;
            8'd137: cosine_value = -125;
            8'd138: cosine_value = -124;
            8'd139: cosine_value = -123;
            8'd140: cosine_value = -122;
            8'd141: cosine_value = -122;
            8'd142: cosine_value = -121;
            8'd143: cosine_value = -119;
            8'd144: cosine_value = -118;
            8'd145: cosine_value = -117;
            8'd146: cosine_value = -116;
            8'd147: cosine_value = -114;
            8'd148: cosine_value = -113;
            8'd149: cosine_value = -111;
            8'd150: cosine_value = -110;
            8'd151: cosine_value = -108;
            8'd152: cosine_value = -106;
            8'd153: cosine_value = -105;
            8'd154: cosine_value = -103;
            8'd155: cosine_value = -101;
            8'd156: cosine_value = -99;
            8'd157: cosine_value = -97;
            8'd158: cosine_value = -95;
            8'd159: cosine_value = -93;
            8'd160: cosine_value = -91;
            8'd161: cosine_value = -88;
            8'd162: cosine_value = -86;
            8'd163: cosine_value = -84;
            8'd164: cosine_value = -81;
            8'd165: cosine_value = -79;
            8'd166: cosine_value = -76;
            8'd167: cosine_value = -74;
            8'd168: cosine_value = -71;
            8'd169: cosine_value = -68;
            8'd170: cosine_value = -66;
            8'd171: cosine_value = -63;
            8'd172: cosine_value = -60;
            8'd173: cosine_value = -58;
            8'd174: cosine_value = -55;
            8'd175: cosine_value = -52;
            8'd176: cosine_value = -49;
            8'd177: cosine_value = -46;
            8'd178: cosine_value = -43;
            8'd179: cosine_value = -40;
            8'd180: cosine_value = -37;
            8'd181: cosine_value = -34;
            8'd182: cosine_value = -31;
            8'd183: cosine_value = -28;
            8'd184: cosine_value = -25;
            8'd185: cosine_value = -22;
            8'd186: cosine_value = -19;
            8'd187: cosine_value = -16;
            8'd188: cosine_value = -13;
            8'd189: cosine_value = -9;
            8'd190: cosine_value = -6;
            8'd191: cosine_value = -3;
            8'd192: cosine_value = 0;
            8'd193: cosine_value = 3;
            8'd194: cosine_value = 6;
            8'd195: cosine_value = 9;
            8'd196: cosine_value = 13;
            8'd197: cosine_value = 16;
            8'd198: cosine_value = 19;
            8'd199: cosine_value = 22;
            8'd200: cosine_value = 25;
            8'd201: cosine_value = 28;
            8'd202: cosine_value = 31;
            8'd203: cosine_value = 34;
            8'd204: cosine_value = 37;
            8'd205: cosine_value = 40;
            8'd206: cosine_value = 43;
            8'd207: cosine_value = 46;
            8'd208: cosine_value = 49;
            8'd209: cosine_value = 52;
            8'd210: cosine_value = 55;
            8'd211: cosine_value = 58;
            8'd212: cosine_value = 60;
            8'd213: cosine_value = 63;
            8'd214: cosine_value = 66;
            8'd215: cosine_value = 68;
            8'd216: cosine_value = 71;
            8'd217: cosine_value = 74;
            8'd218: cosine_value = 76;
            8'd219: cosine_value = 79;
            8'd220: cosine_value = 81;
            8'd221: cosine_value = 84;
            8'd222: cosine_value = 86;
            8'd223: cosine_value = 88;
            8'd224: cosine_value = 91;
            8'd225: cosine_value = 93;
            8'd226: cosine_value = 95;
            8'd227: cosine_value = 97;
            8'd228: cosine_value = 99;
            8'd229: cosine_value = 101;
            8'd230: cosine_value = 103;
            8'd231: cosine_value = 105;
            8'd232: cosine_value = 106;
            8'd233: cosine_value = 108;
            8'd234: cosine_value = 110;
            8'd235: cosine_value = 111;
            8'd236: cosine_value = 113;
            8'd237: cosine_value = 114;
            8'd238: cosine_value = 116;
            8'd239: cosine_value = 117;
            8'd240: cosine_value = 118;
            8'd241: cosine_value = 119;
            8'd242: cosine_value = 121;
            8'd243: cosine_value = 122;
            8'd244: cosine_value = 122;
            8'd245: cosine_value = 123;
            8'd246: cosine_value = 124;
            8'd247: cosine_value = 125;
            8'd248: cosine_value = 126;
            8'd249: cosine_value = 126;
            8'd250: cosine_value = 127;
            8'd251: cosine_value = 127;
            8'd252: cosine_value = 127;
            8'd253: cosine_value = 127;
            8'd254: cosine_value = 127;
            8'd255: cosine_value = 127;
            //default: cosine_value = /* default action */;
        endcase
    end



    






endmodule
